module xnor1(a,b,c);
input a,b;
output c;
xnor(c,a,b);
endmodule