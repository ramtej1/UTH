`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.10.2023 12:39:14
// Design Name: 
// Module Name: Keccak_absorb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Keccak_absorb(string1
    );
    output string1;
reg [63:0]a00=0,a01=0,a02=0,a03=0,a04=0;
reg [63:0]a10=0,a11=0,a12=0,a13=0,a14=0;
reg [63:0]a20=0,a21=0,a22=0,a23=0,a24=0;
reg [63:0]a30=0,a31=0,a32=0,a33=0,a34=0;
reg [63:0]a40=0,a41=0,a42=0,a43=0,a44=0;




endmodule
